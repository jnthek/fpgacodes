module uart 
#(
    parameter DELAY_UNITS = 234
)
(
    input clk,
    output uart_tx,
    input enable_tx
);



endmodule